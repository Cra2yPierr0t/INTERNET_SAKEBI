module internet_sakebi_top (
  input         i_rstn,

  // RMII PHY interface
  input         i_rmii_txclk,
  input  [1:0]  i_rmii_rxd,
  input         i_rmii_crs_dv,
  output [1:0]  o_rmii_txd,
  output        o_rmii_txen
);

  

endmodule
