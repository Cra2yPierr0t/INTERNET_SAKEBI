module internet_sakebi_top_tb;
endmodule
