module internet_sakebi_top (

);
endmodule
